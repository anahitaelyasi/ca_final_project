module datapath(
    input [3:0] R1, R2,
    input E, clk, rst,
    input B1, B2,
    output [3:0] outr 
);


endmodule